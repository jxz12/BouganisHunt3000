module LowC (clk, out);
	input clk;
	output out;
	
reg[14:0] clkDivider = 11;
reg[14:0] counter;

always @(posedge clk)
	if(counter == clkDivider)
		counter <= 1;
	else counter <= counter + 1;
	
reg out;
always @(posedge clk)
	if(counter == 1)
		out <= ~out;

endmodule