module Splitter24 (in, out);
	input in;
	output[23:0] out;

assign out[0] = in;
assign out[1] = in;
assign out[2] = in;
assign out[3] = in;
assign out[4] = in;
assign out[5] = in;
assign out[6] = in;
assign out[7] = in;
assign out[8] = in;
assign out[9] = in;
assign out[10] = in;
assign out[11] = in;
assign out[12] = in;
assign out[13] = in;
assign out[14] = in;
assign out[15] = in;
assign out[16] = in;
assign out[17] = in;
assign out[18] = in;
assign out[19] = in;
assign out[20] = in;
assign out[21] = in;
assign out[22] = in;
assign out[23] = in;

endmodule