module splitter6 (in, out);
	input in;
	output[5:0] out;

assign out[0] = in;
assign out[1] = in;
assign out[2] = in;
assign out[3] = in;
assign out[4] = in;
assign out[5] = in;

endmodule