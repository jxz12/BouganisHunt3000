module eightbitDemux (select, out);
	input [2:0] select;
	output [7:0] out;

assign out[0] = ~select[2] & ~select[1] & ~select[0];
assign out[1] = ~select[2] & ~select[1] & select[0];
assign out[2] = ~select[2] & select[1] & ~select[0];
assign out[3] = ~select[2] & select[1] & select[0];
assign out[4] = select[2] & ~select[1] & ~select[0];
assign out[5] = select[2] & ~select[1] & select[0];
assign out[6] = select[2] & select[1] & ~select[0];
assign out[7] = select[2] & select[1] & select[0];

endmodule