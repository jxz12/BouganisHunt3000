module Splitter (in, out);
	input in;
	output[9:0] out;

assign out[0] = in;
assign out[1] = in;
assign out[2] = in;
assign out[3] = in;
assign out[4] = in;
assign out[5] = in;
assign out[6] = in;
assign out[7] = in;
assign out[8] = in;
assign out[9] = in;

endmodule